`default_nettype none

module log_lut_rom #(
    parameter NUM_SEGMENTS = 64,
    parameter U_WID = 6,
    parameter X_WID = 16
)(
    input wire clk,
    input wire [U_WID-1:0] u_i,
    output bit signed [X_WID-1:0] x_o
);

        always @(posedge clk) begin
        case (u_i)
            (U_WID)'('b000000) : x_o = (X_WID)'('b1001101101000010);
            (U_WID)'('b000001) : x_o = (X_WID)'('b0111100000011011);
            (U_WID)'('b000010) : x_o = (X_WID)'('b0110011111000011);
            (U_WID)'('b000011) : x_o = (X_WID)'('b0101110011111110);
            (U_WID)'('b000100) : x_o = (X_WID)'('b0101010011110100);
            (U_WID)'('b000101) : x_o = (X_WID)'('b0100111010001000);
            (U_WID)'('b000110) : x_o = (X_WID)'('b0100100100101111);
            (U_WID)'('b000111) : x_o = (X_WID)'('b0100010010011011);
            (U_WID)'('b001000) : x_o = (X_WID)'('b0100000010011010);
            (U_WID)'('b001001) : x_o = (X_WID)'('b0011110100001010);
            (U_WID)'('b001010) : x_o = (X_WID)'('b0011100111010111);
            (U_WID)'('b001011) : x_o = (X_WID)'('b0011011011101101);
            (U_WID)'('b001100) : x_o = (X_WID)'('b0011010001000010);
            (U_WID)'('b001101) : x_o = (X_WID)'('b0011000111001100);
            (U_WID)'('b001110) : x_o = (X_WID)'('b0010111110000010);
            (U_WID)'('b001111) : x_o = (X_WID)'('b0010110101100000);
            (U_WID)'('b010000) : x_o = (X_WID)'('b0010101101100000);
            (U_WID)'('b010001) : x_o = (X_WID)'('b0010100101111110);
            (U_WID)'('b010010) : x_o = (X_WID)'('b0010011110110111);
            (U_WID)'('b010011) : x_o = (X_WID)'('b0010011000000111);
            (U_WID)'('b010100) : x_o = (X_WID)'('b0010010001101110);
            (U_WID)'('b010101) : x_o = (X_WID)'('b0010001011101000);
            (U_WID)'('b010110) : x_o = (X_WID)'('b0010000101110011);
            (U_WID)'('b010111) : x_o = (X_WID)'('b0010000000001111);
            (U_WID)'('b011000) : x_o = (X_WID)'('b0001111010111010);
            (U_WID)'('b011001) : x_o = (X_WID)'('b0001110101110010);
            (U_WID)'('b011010) : x_o = (X_WID)'('b0001110000110111);
            (U_WID)'('b011011) : x_o = (X_WID)'('b0001101100000111);
            (U_WID)'('b011100) : x_o = (X_WID)'('b0001100111100011);
            (U_WID)'('b011101) : x_o = (X_WID)'('b0001100011001000);
            (U_WID)'('b011110) : x_o = (X_WID)'('b0001011110110111);
            (U_WID)'('b011111) : x_o = (X_WID)'('b0001011010101111);
            (U_WID)'('b100000) : x_o = (X_WID)'('b0001010110101111);
            (U_WID)'('b100001) : x_o = (X_WID)'('b0001010010110110);
            (U_WID)'('b100010) : x_o = (X_WID)'('b0001001111000110);
            (U_WID)'('b100011) : x_o = (X_WID)'('b0001001011011011);
            (U_WID)'('b100100) : x_o = (X_WID)'('b0001000111111000);
            (U_WID)'('b100101) : x_o = (X_WID)'('b0001000100011010);
            (U_WID)'('b100110) : x_o = (X_WID)'('b0001000001000011);
            (U_WID)'('b100111) : x_o = (X_WID)'('b0000111101110001);
            (U_WID)'('b101000) : x_o = (X_WID)'('b0000111010100100);
            (U_WID)'('b101001) : x_o = (X_WID)'('b0000110111011100);
            (U_WID)'('b101010) : x_o = (X_WID)'('b0000110100011001);
            (U_WID)'('b101011) : x_o = (X_WID)'('b0000110001011011);
            (U_WID)'('b101100) : x_o = (X_WID)'('b0000101110100000);
            (U_WID)'('b101101) : x_o = (X_WID)'('b0000101011101010);
            (U_WID)'('b101110) : x_o = (X_WID)'('b0000101000111000);
            (U_WID)'('b101111) : x_o = (X_WID)'('b0000100110001010);
            (U_WID)'('b110000) : x_o = (X_WID)'('b0000100011011111);
            (U_WID)'('b110001) : x_o = (X_WID)'('b0000100000111000);
            (U_WID)'('b110010) : x_o = (X_WID)'('b0000011110010100);
            (U_WID)'('b110011) : x_o = (X_WID)'('b0000011011110100);
            (U_WID)'('b110100) : x_o = (X_WID)'('b0000011001010110);
            (U_WID)'('b110101) : x_o = (X_WID)'('b0000010110111100);
            (U_WID)'('b110110) : x_o = (X_WID)'('b0000010100100100);
            (U_WID)'('b110111) : x_o = (X_WID)'('b0000010010001111);
            (U_WID)'('b111000) : x_o = (X_WID)'('b0000001111111101);
            (U_WID)'('b111001) : x_o = (X_WID)'('b0000001101101101);
            (U_WID)'('b111010) : x_o = (X_WID)'('b0000001011100000);
            (U_WID)'('b111011) : x_o = (X_WID)'('b0000001001010101);
            (U_WID)'('b111100) : x_o = (X_WID)'('b0000000111001100);
            (U_WID)'('b111101) : x_o = (X_WID)'('b0000000101000110);
            (U_WID)'('b111110) : x_o = (X_WID)'('b0000000011000010);
            (U_WID)'('b111111) : x_o = (X_WID)'('b0000000001000000);
            default: x_o = 0;
        endcase
    end




endmodule: log_lut_rom